LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Count2Cycle IS
   PORT(
			clk           	 	:  IN    STD_LOGIC;                                
			reset          	:  IN    STD_LOGIC; 
			Counter        	:  IN    STD_LOGIC_VECTOR(9 DOWNTO 0);                           
			DutyCycle       	:  OUT   STD_LOGIC_VECTOR(9 DOWNTO 0)
		);  
END Count2Cycle;

ARCHITECTURE behavior OF Count2Cycle IS
	type array_1d is array (0 to 1023) of integer;
	constant C2C_LUT : array_1d := (
(	511	)	,
(	514	)	,
(	517	)	,
(	520	)	,
(	524	)	,
(	527	)	,
(	530	)	,
(	533	)	,
(	536	)	,
(	539	)	,
(	542	)	,
(	545	)	,
(	549	)	,
(	552	)	,
(	555	)	,
(	558	)	,
(	561	)	,
(	564	)	,
(	567	)	,
(	570	)	,
(	574	)	,
(	577	)	,
(	580	)	,
(	583	)	,
(	586	)	,
(	589	)	,
(	592	)	,
(	595	)	,
(	598	)	,
(	602	)	,
(	605	)	,
(	608	)	,
(	611	)	,
(	614	)	,
(	617	)	,
(	620	)	,
(	623	)	,
(	626	)	,
(	629	)	,
(	632	)	,
(	635	)	,
(	638	)	,
(	641	)	,
(	644	)	,
(	647	)	,
(	650	)	,
(	653	)	,
(	656	)	,
(	659	)	,
(	662	)	,
(	665	)	,
(	668	)	,
(	671	)	,
(	674	)	,
(	677	)	,
(	680	)	,
(	683	)	,
(	686	)	,
(	689	)	,
(	692	)	,
(	695	)	,
(	698	)	,
(	701	)	,
(	704	)	,
(	707	)	,
(	710	)	,
(	713	)	,
(	715	)	,
(	718	)	,
(	721	)	,
(	724	)	,
(	727	)	,
(	730	)	,
(	733	)	,
(	735	)	,
(	738	)	,
(	741	)	,
(	744	)	,
(	747	)	,
(	749	)	,
(	752	)	,
(	755	)	,
(	758	)	,
(	760	)	,
(	763	)	,
(	766	)	,
(	769	)	,
(	771	)	,
(	774	)	,
(	777	)	,
(	779	)	,
(	782	)	,
(	785	)	,
(	787	)	,
(	790	)	,
(	793	)	,
(	795	)	,
(	798	)	,
(	800	)	,
(	803	)	,
(	805	)	,
(	808	)	,
(	811	)	,
(	813	)	,
(	816	)	,
(	818	)	,
(	821	)	,
(	823	)	,
(	826	)	,
(	828	)	,
(	831	)	,
(	833	)	,
(	835	)	,
(	838	)	,
(	840	)	,
(	843	)	,
(	845	)	,
(	847	)	,
(	850	)	,
(	852	)	,
(	854	)	,
(	857	)	,
(	859	)	,
(	861	)	,
(	864	)	,
(	866	)	,
(	868	)	,
(	870	)	,
(	873	)	,
(	875	)	,
(	877	)	,
(	879	)	,
(	881	)	,
(	884	)	,
(	886	)	,
(	888	)	,
(	890	)	,
(	892	)	,
(	894	)	,
(	896	)	,
(	898	)	,
(	900	)	,
(	902	)	,
(	904	)	,
(	906	)	,
(	908	)	,
(	910	)	,
(	912	)	,
(	914	)	,
(	916	)	,
(	918	)	,
(	920	)	,
(	922	)	,
(	924	)	,
(	925	)	,
(	927	)	,
(	929	)	,
(	931	)	,
(	933	)	,
(	934	)	,
(	936	)	,
(	938	)	,
(	940	)	,
(	941	)	,
(	943	)	,
(	945	)	,
(	946	)	,
(	948	)	,
(	950	)	,
(	951	)	,
(	953	)	,
(	954	)	,
(	956	)	,
(	957	)	,
(	959	)	,
(	960	)	,
(	962	)	,
(	963	)	,
(	965	)	,
(	966	)	,
(	968	)	,
(	969	)	,
(	970	)	,
(	972	)	,
(	973	)	,
(	975	)	,
(	976	)	,
(	977	)	,
(	978	)	,
(	980	)	,
(	981	)	,
(	982	)	,
(	983	)	,
(	985	)	,
(	986	)	,
(	987	)	,
(	988	)	,
(	989	)	,
(	990	)	,
(	991	)	,
(	992	)	,
(	993	)	,
(	994	)	,
(	995	)	,
(	996	)	,
(	997	)	,
(	998	)	,
(	999	)	,
(	1000	)	,
(	1001	)	,
(	1002	)	,
(	1003	)	,
(	1004	)	,
(	1004	)	,
(	1005	)	,
(	1006	)	,
(	1007	)	,
(	1008	)	,
(	1008	)	,
(	1009	)	,
(	1010	)	,
(	1010	)	,
(	1011	)	,
(	1012	)	,
(	1012	)	,
(	1013	)	,
(	1013	)	,
(	1014	)	,
(	1015	)	,
(	1015	)	,
(	1016	)	,
(	1016	)	,
(	1017	)	,
(	1017	)	,
(	1017	)	,
(	1018	)	,
(	1018	)	,
(	1019	)	,
(	1019	)	,
(	1019	)	,
(	1020	)	,
(	1020	)	,
(	1020	)	,
(	1020	)	,
(	1021	)	,
(	1021	)	,
(	1021	)	,
(	1021	)	,
(	1021	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1022	)	,
(	1021	)	,
(	1021	)	,
(	1021	)	,
(	1021	)	,
(	1021	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1019	)	,
(	1019	)	,
(	1018	)	,
(	1018	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1016	)	,
(	1015	)	,
(	1015	)	,
(	1014	)	,
(	1014	)	,
(	1013	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	971	)	,
(	970	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	964	)	,
(	963	)	,
(	961	)	,
(	960	)	,
(	958	)	,
(	957	)	,
(	955	)	,
(	954	)	,
(	952	)	,
(	950	)	,
(	949	)	,
(	947	)	,
(	946	)	,
(	944	)	,
(	942	)	,
(	940	)	,
(	939	)	,
(	937	)	,
(	935	)	,
(	934	)	,
(	932	)	,
(	930	)	,
(	928	)	,
(	926	)	,
(	925	)	,
(	923	)	,
(	921	)	,
(	919	)	,
(	917	)	,
(	915	)	,
(	913	)	,
(	911	)	,
(	909	)	,
(	907	)	,
(	905	)	,
(	903	)	,
(	901	)	,
(	899	)	,
(	897	)	,
(	895	)	,
(	893	)	,
(	891	)	,
(	889	)	,
(	887	)	,
(	885	)	,
(	882	)	,
(	880	)	,
(	878	)	,
(	876	)	,
(	874	)	,
(	872	)	,
(	869	)	,
(	867	)	,
(	865	)	,
(	863	)	,
(	860	)	,
(	858	)	,
(	856	)	,
(	853	)	,
(	851	)	,
(	849	)	,
(	846	)	,
(	844	)	,
(	841	)	,
(	839	)	,
(	837	)	,
(	834	)	,
(	832	)	,
(	829	)	,
(	827	)	,
(	824	)	,
(	822	)	,
(	819	)	,
(	817	)	,
(	814	)	,
(	812	)	,
(	809	)	,
(	807	)	,
(	804	)	,
(	802	)	,
(	799	)	,
(	796	)	,
(	794	)	,
(	791	)	,
(	789	)	,
(	786	)	,
(	783	)	,
(	781	)	,
(	778	)	,
(	775	)	,
(	773	)	,
(	770	)	,
(	767	)	,
(	764	)	,
(	762	)	,
(	759	)	,
(	756	)	,
(	754	)	,
(	751	)	,
(	748	)	,
(	745	)	,
(	742	)	,
(	740	)	,
(	737	)	,
(	734	)	,
(	731	)	,
(	728	)	,
(	725	)	,
(	723	)	,
(	720	)	,
(	717	)	,
(	714	)	,
(	711	)	,
(	708	)	,
(	705	)	,
(	702	)	,
(	700	)	,
(	697	)	,
(	694	)	,
(	691	)	,
(	688	)	,
(	685	)	,
(	682	)	,
(	679	)	,
(	676	)	,
(	673	)	,
(	670	)	,
(	667	)	,
(	664	)	,
(	661	)	,
(	658	)	,
(	655	)	,
(	652	)	,
(	649	)	,
(	646	)	,
(	643	)	,
(	640	)	,
(	637	)	,
(	634	)	,
(	631	)	,
(	628	)	,
(	625	)	,
(	622	)	,
(	619	)	,
(	615	)	,
(	612	)	,
(	609	)	,
(	606	)	,
(	603	)	,
(	600	)	,
(	597	)	,
(	594	)	,
(	591	)	,
(	588	)	,
(	585	)	,
(	581	)	,
(	578	)	,
(	575	)	,
(	572	)	,
(	569	)	,
(	566	)	,
(	563	)	,
(	560	)	,
(	556	)	,
(	553	)	,
(	550	)	,
(	547	)	,
(	544	)	,
(	541	)	,
(	538	)	,
(	535	)	,
(	531	)	,
(	528	)	,
(	525	)	,
(	522	)	,
(	519	)	,
(	516	)	,
(	513	)	,
(	509	)	,
(	506	)	,
(	503	)	,
(	500	)	,
(	497	)	,
(	494	)	,
(	491	)	,
(	488	)	,
(	484	)	,
(	481	)	,
(	478	)	,
(	475	)	,
(	472	)	,
(	469	)	,
(	466	)	,
(	462	)	,
(	459	)	,
(	456	)	,
(	453	)	,
(	450	)	,
(	447	)	,
(	444	)	,
(	441	)	,
(	438	)	,
(	434	)	,
(	431	)	,
(	428	)	,
(	425	)	,
(	422	)	,
(	419	)	,
(	416	)	,
(	413	)	,
(	410	)	,
(	407	)	,
(	404	)	,
(	401	)	,
(	397	)	,
(	394	)	,
(	391	)	,
(	388	)	,
(	385	)	,
(	382	)	,
(	379	)	,
(	376	)	,
(	373	)	,
(	370	)	,
(	367	)	,
(	364	)	,
(	361	)	,
(	358	)	,
(	355	)	,
(	352	)	,
(	349	)	,
(	346	)	,
(	343	)	,
(	340	)	,
(	337	)	,
(	334	)	,
(	331	)	,
(	328	)	,
(	326	)	,
(	323	)	,
(	320	)	,
(	317	)	,
(	314	)	,
(	311	)	,
(	308	)	,
(	305	)	,
(	302	)	,
(	299	)	,
(	297	)	,
(	294	)	,
(	291	)	,
(	288	)	,
(	285	)	,
(	282	)	,
(	280	)	,
(	277	)	,
(	274	)	,
(	271	)	,
(	269	)	,
(	266	)	,
(	263	)	,
(	260	)	,
(	258	)	,
(	255	)	,
(	252	)	,
(	249	)	,
(	247	)	,
(	244	)	,
(	241	)	,
(	239	)	,
(	236	)	,
(	233	)	,
(	231	)	,
(	228	)	,
(	226	)	,
(	223	)	,
(	220	)	,
(	218	)	,
(	215	)	,
(	213	)	,
(	210	)	,
(	208	)	,
(	205	)	,
(	203	)	,
(	200	)	,
(	198	)	,
(	195	)	,
(	193	)	,
(	190	)	,
(	188	)	,
(	185	)	,
(	183	)	,
(	181	)	,
(	178	)	,
(	176	)	,
(	173	)	,
(	171	)	,
(	169	)	,
(	166	)	,
(	164	)	,
(	162	)	,
(	160	)	,
(	157	)	,
(	155	)	,
(	153	)	,
(	151	)	,
(	148	)	,
(	146	)	,
(	144	)	,
(	142	)	,
(	140	)	,
(	137	)	,
(	135	)	,
(	133	)	,
(	131	)	,
(	129	)	,
(	127	)	,
(	125	)	,
(	123	)	,
(	121	)	,
(	119	)	,
(	117	)	,
(	115	)	,
(	113	)	,
(	111	)	,
(	109	)	,
(	107	)	,
(	105	)	,
(	103	)	,
(	101	)	,
(	99	)	,
(	98	)	,
(	96	)	,
(	94	)	,
(	92	)	,
(	90	)	,
(	89	)	,
(	87	)	,
(	85	)	,
(	83	)	,
(	82	)	,
(	80	)	,
(	78	)	,
(	77	)	,
(	75	)	,
(	73	)	,
(	72	)	,
(	70	)	,
(	68	)	,
(	67	)	,
(	65	)	,
(	64	)	,
(	62	)	,
(	61	)	,
(	59	)	,
(	58	)	,
(	56	)	,
(	55	)	,
(	54	)	,
(	52	)	,
(	51	)	,
(	50	)	,
(	48	)	,
(	47	)	,
(	46	)	,
(	44	)	,
(	43	)	,
(	42	)	,
(	41	)	,
(	39	)	,
(	38	)	,
(	37	)	,
(	36	)	,
(	35	)	,
(	33	)	,
(	32	)	,
(	31	)	,
(	30	)	,
(	29	)	,
(	28	)	,
(	27	)	,
(	26	)	,
(	25	)	,
(	24	)	,
(	23	)	,
(	22	)	,
(	21	)	,
(	20	)	,
(	20	)	,
(	19	)	,
(	18	)	,
(	17	)	,
(	16	)	,
(	16	)	,
(	15	)	,
(	14	)	,
(	13	)	,
(	13	)	,
(	12	)	,
(	11	)	,
(	11	)	,
(	10	)	,
(	9	)	,
(	9	)	,
(	8	)	,
(	8	)	,
(	7	)	,
(	7	)	,
(	6	)	,
(	6	)	,
(	5	)	,
(	5	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	4	)	,
(	4	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	6	)	,
(	6	)	,
(	7	)	,
(	7	)	,
(	8	)	,
(	8	)	,
(	9	)	,
(	10	)	,
(	10	)	,
(	11	)	,
(	12	)	,
(	12	)	,
(	13	)	,
(	14	)	,
(	14	)	,
(	15	)	,
(	16	)	,
(	17	)	,
(	17	)	,
(	18	)	,
(	19	)	,
(	20	)	,
(	21	)	,
(	22	)	,
(	23	)	,
(	24	)	,
(	25	)	,
(	26	)	,
(	27	)	,
(	28	)	,
(	29	)	,
(	30	)	,
(	31	)	,
(	32	)	,
(	33	)	,
(	34	)	,
(	35	)	,
(	36	)	,
(	37	)	,
(	39	)	,
(	40	)	,
(	41	)	,
(	42	)	,
(	44	)	,
(	45	)	,
(	46	)	,
(	47	)	,
(	49	)	,
(	50	)	,
(	51	)	,
(	53	)	,
(	54	)	,
(	56	)	,
(	57	)	,
(	59	)	,
(	60	)	,
(	62	)	,
(	63	)	,
(	65	)	,
(	66	)	,
(	68	)	,
(	69	)	,
(	71	)	,
(	72	)	,
(	74	)	,
(	76	)	,
(	77	)	,
(	79	)	,
(	81	)	,
(	82	)	,
(	84	)	,
(	86	)	,
(	88	)	,
(	89	)	,
(	91	)	,
(	93	)	,
(	95	)	,
(	97	)	,
(	98	)	,
(	100	)	,
(	102	)	,
(	104	)	,
(	106	)	,
(	108	)	,
(	110	)	,
(	112	)	,
(	114	)	,
(	116	)	,
(	118	)	,
(	120	)	,
(	122	)	,
(	124	)	,
(	126	)	,
(	128	)	,
(	130	)	,
(	132	)	,
(	134	)	,
(	136	)	,
(	138	)	,
(	141	)	,
(	143	)	,
(	145	)	,
(	147	)	,
(	149	)	,
(	152	)	,
(	154	)	,
(	156	)	,
(	158	)	,
(	161	)	,
(	163	)	,
(	165	)	,
(	167	)	,
(	170	)	,
(	172	)	,
(	175	)	,
(	177	)	,
(	179	)	,
(	182	)	,
(	184	)	,
(	186	)	,
(	189	)	,
(	191	)	,
(	194	)	,
(	196	)	,
(	199	)	,
(	201	)	,
(	204	)	,
(	206	)	,
(	209	)	,
(	211	)	,
(	214	)	,
(	216	)	,
(	219	)	,
(	222	)	,
(	224	)	,
(	227	)	,
(	229	)	,
(	232	)	,
(	235	)	,
(	237	)	,
(	240	)	,
(	243	)	,
(	245	)	,
(	248	)	,
(	251	)	,
(	253	)	,
(	256	)	,
(	259	)	,
(	262	)	,
(	264	)	,
(	267	)	,
(	270	)	,
(	273	)	,
(	275	)	,
(	278	)	,
(	281	)	,
(	284	)	,
(	287	)	,
(	289	)	,
(	292	)	,
(	295	)	,
(	298	)	,
(	301	)	,
(	304	)	,
(	307	)	,
(	309	)	,
(	312	)	,
(	315	)	,
(	318	)	,
(	321	)	,
(	324	)	,
(	327	)	,
(	330	)	,
(	333	)	,
(	336	)	,
(	339	)	,
(	342	)	,
(	345	)	,
(	347	)	,
(	350	)	,
(	353	)	,
(	356	)	,
(	359	)	,
(	362	)	,
(	365	)	,
(	368	)	,
(	371	)	,
(	374	)	,
(	378	)	,
(	381	)	,
(	384	)	,
(	387	)	,
(	390	)	,
(	393	)	,
(	396	)	,
(	399	)	,
(	402	)	,
(	405	)	,
(	408	)	,
(	411	)	,
(	414	)	,
(	417	)	,
(	420	)	,
(	423	)	,
(	427	)	,
(	430	)	,
(	433	)	,
(	436	)	,
(	439	)	,
(	442	)	,
(	445	)	,
(	448	)	,
(	451	)	,
(	455	)	,
(	458	)	,
(	461	)	,
(	464	)	,
(	467	)	,
(	470	)	,
(	473	)	,
(	476	)	,
(	480	)	,
(	483	)	,
(	486	)	,
(	489	)	,
(	492	)	,
(	495	)	,
(	498	)	,
(	501	)	,
(	505	)	,
(	508	)	,
(	511	)	
);
begin
process (clk, reset)
begin
	if rising_edge(clk) then
		if reset = '1' then
			DutyCycle <= (others => '0');
		else
			DutyCycle <= std_logic_vector(to_unsigned(C2C_LUT(to_integer(unsigned(Counter))),DutyCycle'Length));
		end if;
	end if;
end process;
	
	
end behavior;