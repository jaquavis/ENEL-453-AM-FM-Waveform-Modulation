LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Distance2Offset IS
   PORT(
			clk            :  IN    STD_LOGIC;                                
			reset          :  IN    STD_LOGIC; 
			distance       :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
			offset         :  OUT   STD_LOGIC_VECTOR(9 DOWNTO 0)
		  );  
END Distance2Offset;

ARCHITECTURE behavior OF Distance2Offset IS

type array_1d is array (0 to 4095) of integer;

constant D2O_LUT : array_1d := ( 
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	852	)
);
begin

process (clk, reset)
begin
	if rising_edge(clk) then
		if reset = '1' then
			offset <= (others => '0');
		else
			offset <= std_logic_vector(to_unsigned(D2O_LUT(to_integer(unsigned(distance))),offset'length));
		end if;
	end if;
end process;

end behavior;